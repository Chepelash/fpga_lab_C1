module packet_classer_tb;



endmodule
